module driver7seg (b,d);

	input [3:0] b; //número a ser mostrado
	output reg [6:0] d; //saida de 7 segmentos

	always @* begin
	
		case (b)
			
			4'd0: d = 7'b1000000; //0
			4'd1: d = 7'b1111001; //1
			4'd2: d = 7'b0100100; //2
			4'd3: d = 7'b0110000; //3
			4'd4: d = 7'b0011001; //4
			4'd5: d = 7'b0010010; //5
			4'd6: d = 7'b0000010; //6
			4'd7: d = 7'b1111000; //7
			4'd8: d = 7'b0000000; //8
			4'd9: d = 7'b0010000; //9

		endcase
	
	end


endmodule
